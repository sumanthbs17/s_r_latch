interface intf();
    // ------------------- port declaration-------------------------------------
    logic s;
    logic r;
    logic q;
    logic qbar;
    //--------------------------------------------------------------------------
    //--------------------------------------------------------------------------
        
endinterface
